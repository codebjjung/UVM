module UART (
