class sequence_item extends uvm_sequence_item
	`uvm_object_utils(sequence_item)
