class monitor extends
